
module HeaderCreatorN6ToN3(
  input logic             CLK,
  input logic             reset,
  input logic   [31 : 0]  bus,
  output logic  [15 : 0]  bus_read_id, 
  output logic            read_bus_req,           
  input HC_N6_to_N3       hc_fields
);




endmodule