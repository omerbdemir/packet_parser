`define BUS_WIDTH_B         4
`define BYTE_WIDTH          8
`define BUS_WIDTH_BITS      (`BUS_WIDTH_B * `BYTE_WIDTH)
