
module HeaderCreatorN6ToN3(
  input logic CLK,
  input logic reset,
  input HC_N6_to_N3
);



endmodule