module HeaderCreatorN3ToN6(
  input logic CLK,
  input logic reset,
  input HC_N3_to_N6
);

endmodule