package my_package;
  import my_test_lib::*;
endpackage