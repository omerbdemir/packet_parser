module HeaderCreatorN3ToN6(
  input logic CLK,
  input logic reset,
  input logic   [31 : 0]  bus,
  output logic  [15 : 0]  bus_read_id,
  output logic            bus_read_req,
  input HC_N3_to_N6
);

endmodule